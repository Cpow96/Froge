module blogrom
(
	input logic [6:0] DX, DY,
	input logic  dir,
	output logic [7:0] data
);
// 1
	int blog [24][96];
	
	always_ff
	begin
	
	blog = '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,26,26,26,26,26,26,26,26,26,26,26,27,27,27,27,26,26,26,26,26,26,27,27,26,26,26,26,27,27,26,26,26,26,26,26,26,26,26,26,27,27,27,27,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,27,27,27,27,26,26,26,26,26,26,27,27,26,26,26,26,27,27,26,26,26,26,26,26,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,26,26,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,26,26,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,26,26,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,28,28,29,29,0,0,0,0,0,0,0},
'{0,0,0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,29,28,29,29,0,0,0,0,0},
'{0,0,0,26,26,27,27,27,27,27,28,28,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,29,29,29,27,27,29,29,27,27,27,27,28,28,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,29,29,29,27,27,29,29,27,27,27,27,27,29,27,28,28,27,29,0,0,0,0},
'{0,0,0,26,26,27,27,28,28,28,28,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,27,27,27,29,29,29,29,27,27,28,28,28,28,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,28,28,28,28,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,27,27,27,29,29,29,29,27,27,27,27,27,29,28,29,29,28,27,29,29,0,0,0},
'{0,0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,29,28,28,28,28,28,27,29,0,0,0},
'{0,0,26,26,27,27,27,27,29,29,29,27,27,27,27,27,27,27,27,27,27,27,29,29,29,29,29,27,27,27,27,27,27,27,27,27,29,29,29,27,26,26,26,26,26,27,27,27,27,27,29,29,29,29,27,29,29,29,27,27,27,27,27,27,27,27,27,27,27,29,29,29,29,29,27,27,27,27,27,27,27,27,27,27,29,28,27,28,27,28,28,27,29,29,0,0},
'{0,0,26,26,27,29,29,29,29,27,27,27,27,27,27,27,27,29,29,29,29,29,29,27,27,27,27,27,28,28,28,28,28,28,28,29,29,27,27,27,27,27,27,27,26,29,29,29,29,29,29,27,27,27,29,29,27,27,27,27,27,27,27,27,29,29,29,29,29,29,27,27,27,27,27,28,28,28,28,28,28,28,27,27,29,28,28,27,29,29,28,27,28,29,0,0},
'{0,0,26,26,27,27,27,27,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,27,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,27,28,29,28,28,27,27,29,28,27,28,29,0,0},
'{0,0,26,26,27,27,27,27,27,27,27,27,28,28,28,28,27,27,27,27,27,27,28,28,28,27,27,26,26,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,27,27,27,27,27,27,28,28,28,27,27,27,27,27,27,28,28,28,28,27,27,27,27,27,27,28,28,28,27,27,26,26,27,27,27,27,27,27,27,27,29,29,28,28,27,29,28,28,28,29,0,0},
'{0,0,26,26,26,26,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,27,27,27,27,26,26,26,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,27,27,27,27,26,26,26,27,27,27,27,29,29,27,28,28,27,28,28,27,29,29,0,0},
'{0,0,26,26,27,26,26,26,26,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,29,27,27,27,28,26,26,29,0,0,0},
'{0,0,26,26,27,27,26,26,27,27,26,27,27,27,27,27,27,27,27,27,29,29,27,27,27,27,27,27,27,28,28,28,28,28,27,27,27,26,26,26,27,27,27,27,27,27,26,26,29,29,27,27,27,27,27,27,27,27,26,26,27,27,27,27,27,27,26,29,29,27,27,27,27,27,27,27,28,28,28,28,28,27,27,29,29,27,27,27,28,28,27,26,29,0,0,0},
'{0,0,26,26,27,27,27,27,27,29,29,29,27,27,27,27,27,27,27,29,29,29,29,29,27,27,27,27,27,27,27,27,27,28,28,27,27,29,29,26,26,26,26,26,26,26,26,29,29,29,29,29,27,27,27,27,29,29,29,26,26,26,26,26,26,26,26,29,29,29,29,27,27,27,27,27,27,27,27,27,28,28,27,29,27,27,28,27,28,26,27,26,29,0,0,0},
'{0,0,26,26,27,27,27,27,27,27,27,27,29,29,29,29,29,29,29,29,27,27,27,29,29,27,27,27,27,27,27,27,27,27,28,27,27,27,27,27,29,29,29,29,29,29,29,29,27,27,27,29,29,27,27,27,27,27,27,29,29,29,29,29,29,29,29,27,27,27,29,29,27,27,27,27,27,27,27,27,27,28,2,29,27,27,28,28,28,27,26,29,29,0,0,0},
'{0,0,26,26,27,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,27,27,27,27,27,28,28,27,27,27,27,27,26,26,26,26,26,27,27,27,27,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,27,27,27,27,27,27,29,29,27,27,28,27,26,26,29,0,0,0,0},
'{0,0,0,26,27,27,26,26,28,28,27,27,27,27,27,27,27,27,27,27,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,26,28,28,27,27,27,27,27,27,27,27,27,27,28,28,28,27,27,27,26,28,28,27,27,27,27,27,27,27,27,27,27,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,28,28,29,26,26,29,29,0,0,0,0},
'{0,0,0,26,26,27,27,27,27,27,28,28,28,28,28,28,28,28,28,28,27,27,27,27,27,27,27,26,26,26,26,27,27,27,27,27,27,27,28,28,28,28,28,28,28,28,28,28,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,28,28,28,27,27,27,27,27,27,27,26,26,26,26,27,27,27,27,27,27,29,28,28,26,29,29,0,0,0,0,0,0},
'{0,0,0,26,26,26,26,27,27,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,27,27,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,27,27,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,29,29,29,29,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};

	end
	
	always_ff
	begin
		data = blog[DY][DX];
	//unique case (dir)
		//1'd0: data = truckleft[DY][DX];
		//1'd1: data = truckright[DY][DX];
		
	//endcase

	end
endmodule
