module pacmanJr_ROM
(
	input logic [4:0] addr,
	output logic [31:0] data
);
// 1
	parameter [0:31][31:0] pacROM = {32'b00000000000000000000000000000000,
												32'b00000000000000000000000000000000,
												32'b00000000001111111111110000000000,
												32'b00000000001111111111110000000000,
												32'b00000011111111111111111111000000,
												32'b00000011111111111111111111000000,
												32'b00001111111111111111111111110000,
												32'b00001111111111111111111111110000,
												32'b00111111111111111111111111111100,
												32'b00111111111111111111111111111100,
												32'b11111111111111111111111111111100,
												32'b11111111111111111111111111111100,
												32'b11111111111111111111110000000000,
												32'b11111111111111111111110000000000,
												32'b11111111111111000000000000000000,
												32'b11111111111111000000000000000000,
												32'b11111111111111000000000000000000,
												32'b11111111111111000000000000000000,
												32'b11111111111111111111110000000000,
												32'b11111111111111111111110000000000,
												32'b11111111111111111111111111111100,
												32'b11111111111111111111111111111100,
												32'b00111111111111111111111111111100,
												32'b00111111111111111111111111111100,
												32'b00001111111111111111111111110000,
												32'b00001111111111111111111111110000,
												32'b00000011111111111111111111000000,
												32'b00000011111111111111111111000000,
												32'b00000000001111111111110000000000,
												32'b00000000001111111111110000000000,
												32'b00000000000000000000000000000000,
												32'b00000000000000000000000000000000};

	assign data = pacROM[addr];
												
endmodule
