module slogrom
(
	input logic [5:0] DX, DY,
	input logic  dir,
	output logic [7:0] data
);
// 1
	int slog [24][48];
	
	always_ff
	begin
	
	slog = '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,26,26,26,26,26,26,26,26,26,26,26,27,27,27,27,26,26,26,26,26,26,27,27,26,26,26,26,27,27,26,26,26,26,26,26,0,0,0,0,0,0,0,0},
'{0,0,0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,26,26,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,28,28,29,29,0,0,0,0,0,0},
'{0,0,0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,29,2,29,29,0,0,0,0},
'{0,0,0,26,26,27,27,27,27,27,28,28,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,29,29,29,27,27,29,29,27,27,27,27,27,29,27,28,28,27,29,0,0,0},
'{0,0,0,26,26,27,27,28,28,28,28,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,27,27,27,29,29,29,29,27,27,27,27,27,29,2,29,29,28,27,29,29,0,0},
'{0,0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,29,28,28,28,28,2,27,29,0,0},
'{0,0,26,26,27,27,27,27,29,29,29,27,27,27,27,27,27,27,27,27,27,27,29,29,29,29,29,27,27,27,27,27,27,27,27,27,27,29,2,27,28,27,28,28,27,29,0,0},
'{0,0,26,26,27,29,29,29,29,27,27,27,27,27,27,27,27,29,29,29,29,29,29,27,27,27,27,27,28,28,28,28,28,28,28,27,27,29,28,28,27,29,2,28,27,2,29,0},
'{0,0,26,26,27,27,27,27,28,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,27,28,29,28,28,27,27,29,28,27,28,29,0},
'{0,0,26,26,27,27,27,27,27,27,27,27,28,28,28,28,27,27,27,27,27,27,28,28,28,27,27,26,26,27,27,27,27,27,27,27,27,2,29,28,28,27,29,28,28,28,2,0},
'{0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,28,27,27,27,27,27,27,26,26,26,27,27,27,27,27,29,27,28,28,27,28,28,27,29,29,0},
'{0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,2,29,27,27,27,28,26,26,29,0,0},
'{0,0,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,29,27,27,27,27,27,27,27,28,28,28,28,28,27,27,29,29,27,27,27,28,28,27,26,29,0,0},
'{0,0,26,26,27,27,27,27,27,29,29,29,27,27,27,27,27,27,27,29,29,29,29,29,27,27,27,27,27,27,27,27,27,28,28,27,29,27,27,28,27,28,26,27,26,2,0,0},
'{0,0,26,26,27,27,27,27,27,27,27,27,29,29,29,29,29,29,29,29,27,27,27,29,29,27,27,27,27,27,27,27,27,27,28,2,29,27,27,28,28,28,27,26,2,0,0,0},
'{0,0,26,26,27,28,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,27,27,27,27,27,27,29,29,27,27,28,27,2,26,29,0,0,0},
'{0,0,0,26,27,27,26,26,28,28,27,27,27,27,27,27,27,27,27,27,28,28,28,27,27,27,27,27,27,27,27,27,27,27,27,27,27,29,28,28,29,26,26,29,29,0,0,0},
'{0,0,0,26,26,27,27,27,27,27,28,28,28,28,28,28,28,28,28,28,27,27,27,27,27,27,27,26,26,26,26,27,27,27,27,27,27,2,28,28,26,29,2,29,0,0,0,0},
'{0,0,0,26,26,26,26,27,27,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,29,29,29,2,0,29,29,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};

	end
	
	always_ff
	begin
		data = slog[DY][DX];
	//unique case (dir)
		//1'd0: data = truckleft[DY][DX];
		//1'd1: data = truckright[DY][DX];
		
	//endcase

	end
endmodule
