module map_ROM
(
	input logic [9:0] currX, currY,
	output logic [7:0] outR, outG, outB
);
	// # of map sprites: 20
	// this array holds information on how the map is pieced together from sprites; numbers indicate different sprites of the map
	parameter bit [4:0] map_Layout [0:9][27:0] = '{'{5'd0, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd19, 5'd20, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd2},							// row 0
													 '{5'd3, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd5, 5'd6, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd7},							// row 1
													 '{5'd3, 5'd4, 5'd8, 5'd9, 5'd9, 5'd10, 5'd4, 5'd8, 5'd9, 5'd9, 5'd9, 5'd10, 5'd4, 5'd5, 5'd6, 5'd4, 5'd8, 5'd9, 5'd9, 5'd9, 5'd10, 5'd4, 5'd8, 5'd9, 5'd9, 5'd10, 5'd4, 5'd7},						// row 2
													 '{5'd3, 5'd4, 5'd5, 5'd4, 5'd4, 5'd6, 5'd4, 5'd5, 5'd4, 5'd4, 5'd4, 5'd6, 5'd4, 5'd5, 5'd6, 5'd4, 5'd5, 5'd4, 5'd4, 5'd4, 5'd6, 5'd4, 5'd5, 5'd4, 5'd4, 5'd6, 5'd4, 5'd7},							// row 3
													 '{5'd3, 5'd4, 5'd11, 5'd12, 5'd12, 5'd13, 5'd4, 5'd11, 5'd12, 5'd12, 5'd12, 5'd13, 5'd4, 5'd5, 5'd6, 5'd4, 5'd11, 5'd12, 5'd12, 5'd12, 5'd13, 5'd4, 5'd11, 5'd12, 5'd12, 5'd13, 5'd4, 5'd7},	// row 4
													 '{5'd3, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd7},							// row 5
													 '{5'd3, 5'd4, 5'd8, 5'd9, 5'd9, 5'd10, 5'd4, 5'd8, 5'd10, 5'd4, 5'd8, 5'd9, 5'd9, 5'd9, 5'd9, 5'd9, 5'd9, 5'd10, 5'd4, 5'd8, 5'd10, 5'd4, 5'd8, 5'd9, 5'd9, 5'd10, 5'd4, 5'd7},						// row 6
													 '{5'd3, 5'd4, 5'd11, 5'd12, 5'd12, 5'd13, 5'd4, 5'd5, 5'd6, 5'd4, 5'd11, 5'd12, 5'd12, 5'd10, 5'd8, 5'd12, 5'd12, 5'd13, 5'd4, 5'd5, 5'd6, 5'd4, 5'd11, 5'd12, 5'd12, 5'd13, 5'd4, 5'd7},		// row 7
													 '{5'd3, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd5, 5'd6, 5'd4, 5'd4, 5'd4, 5'd4, 5'd5, 5'd6, 5'd4, 5'd4, 5'd4, 5'd4, 5'd5, 5'd6, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd4, 5'd7},							// row 8
													 '{5'd14, 5'd15, 5'd15, 5'd15, 5'd15, 5'd10, 5'd4, 5'd5, 5'd16, 5'd9, 5'd9, 5'd10, 5'd4, 5'd5, 5'd6, 5'd4, 5'd8, 5'd9, 5'd9, 5'd17, 5'd6, 5'd4, 5'd8, 5'd15, 5'd15, 5'd15, 5'd15, 5'd18}};		// row 9
													 
//	parameter bit [4:0] map_Layout [0:1][27:0] = '{'{5'd0, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd19, 5'd20, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd2},							// row 0
//													 '{5'd0, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd19, 5'd20, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd1, 5'd2}};		// row 9
//													 

		parameter [0:7][7:0] map_0 = {8'b00001111,
											8'b00110000,
											8'b01000000,
											8'b01000111,
											8'b10001000,
											8'b10010000,
											8'b10010000,
											8'b10010000};
//	parameter [0:15][15:0] map_0 = {8'b0000000011111111,
//											8'b0000000011111111,
//											8'b0000111100000000,
//											8'b0000111100000000,
//											8'b0011000000000000,
//											8'b0011000000000000,
//											8'b0011000000111111,
//											8'b0011000000111111,
//											8'b1100000011000000,
//											8'b1100000011000000,
//											8'b1100001100000000,
//											8'b1100001100000000,
//											8'b1100001100000000,
//											8'b1100001100000000,
//											8'b1100001100000000,
//											8'b1100001100000000};
			
	parameter [0:7][7:0] map_1 = {8'b11111111,
											8'b00000000,
											8'b00000000,
											8'b11111111,
											8'b00000000,
											8'b00000000,
											8'b00000000,
											8'b00000000};			
//	parameter [0:15][15:0] map_1 = {8'b1111111111111111,
//											8'b1111111111111111,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b1111111111111111,
//											8'b1111111111111111,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000,
//											8'b0000000000000000};
											
	parameter [0:7][7:0] map_19 = {8'b11111111,
											 8'b00000000,
											 8'b00000000,
											 8'b11000000,
											 8'b00100000,
											 8'b00010000,
											 8'b00010000,
											 8'b00010000};
//	parameter [0:15][15:0] map_19 = {8'b1111111111111111,
//											 8'b1111111111111111,
//											 8'b0000000000000000,
//											 8'b0000000000000000,
//											 8'b0000000000000000,
//											 8'b0000000000000000,
//											 8'b1111000000000000,
//											 8'b1111000000000000,
//											 8'b0000110000000000,
//											 8'b0000110000000000,
//											 8'b0000001100000000,
//											 8'b0000001100000000,
//											 8'b0000001100000000,
//											 8'b0000001100000000,
//											 8'b0000001100000000,
//											 8'b0000001100000000};

	parameter [0:7][7:0] map_20 = {8'b11111111,
											 8'b00000000,
											 8'b00000000,
											 8'b00000011,
											 8'b00000100,
											 8'b00001000,
											 8'b00001000,
											 8'b00001000};

//	parameter [0:15][15:0] map_20 = {8'b1111111111111111,
//											 8'b1111111111111111,
//											 8'b0000000000000000,
//											 8'b0000000000000000,
//											 8'b0000000000000000,
//											 8'b0000000000000000,
//											 8'b0000000000001111,
//											 8'b0000000000001111,
//											 8'b0000000000110000,
//											 8'b0000000000110000,
//											 8'b0000000011000000,
//											 8'b0000000011000000,
//											 8'b0000000011000000,
//											 8'b0000000011000000,
//											 8'b0000000011000000,
//											 8'b0000000011000000};
											 
	parameter [0:7][7:0] map_2 = {8'b11110000,
											8'b00001100,
											8'b00000010,
											8'b11100010,
											8'b00010001,
											8'b00001001,
											8'b00001001,
											8'b00001001};
//	parameter [0:15][15:0] map_2 = {8'b1111111100000000,
//											8'b1111111100000000,
//											8'b0000000011110000,
//											8'b0000000011110000,
//											8'b0000000000001100,
//											8'b0000000000001100,
//											8'b1111110000001100,
//											8'b1111110000001100,
//											8'b0000001100000011,
//											8'b0000001100000011,
//											8'b0000000011000011,
//											8'b0000000011000011,
//											8'b0000000011000011,
//											8'b0000000011000011,
//											8'b0000000011000011,	
//											8'b0000000011000011};	
//										
// 1
//	assign data = mapROM[addr];

	// translate coordinates to a 40x30 grid system
	logic [4:0] indexX, indexY;
	logic [4:0] mapSprite, x, y;
	logic [7:0] spriteData;
	assign y = currY >> 10'd3;
	assign x = currX >> 10'd3;
	assign indexX = currX & 10'd7;//currX % 10'd8;
	assign indexY = currY & 10'd7;//currY % 10'd8;
//	assign indexX = currX % 10'd8;
//	assign indexY = currY % 10'd8;
	assign mapSprite = map_Layout[y][27-x];
//   assign mapSprite = 5'd1;
	
	always_comb begin
	spriteData = 8'd0;
	unique case (mapSprite)
		5'd0: begin
			spriteData = map_0[indexY];
			if (spriteData[7-indexX])
			begin
				// red
				outR = 8'hff;//8'h00;
				outG = 8'h00;
				outB = 8'h00;//8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		5'd1: begin
			spriteData = map_1[indexY];
			if (spriteData[7-indexX])
			begin
				// green
				outR = 8'h00;
				outG = 8'hff;//8'h00;
				outB = 8'h00;//8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		5'd2: begin
			spriteData = map_2[indexY];
			if (spriteData[7-indexX])
			begin
				// yellow
				outR = 8'hff;//8'h00;
				outG = 8'hff;//8'h00;
				outB = 8'h00;//8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		5'd19: begin
			spriteData = map_19[indexY];
			if (spriteData[7-indexX])
			begin
				// orange
				outR = 8'hff;//8'h00;
				outG = 8'ha5;//8'h00;
				outB = 8'h00;//8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		5'd20: begin
			spriteData = map_20[indexY];
			if (spriteData[7-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		default: begin
			outR = 8'hff;
			outG = 8'hff;
			outB = 8'hff;
		end
	endcase
	end
	
endmodule
