module carleftrom
(
	input logic [5:0] DX, DY,
	input logic  dir,
	output logic [7:0] data
);
// 1
	int carleft [24][24];
	
	always_ff
	begin
	
	carleft = '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,6,6,6,6,6,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,6,6,6,0,0,0,6,6,6,6,6,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,6,6,6,0,0,0,0,0,6,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,6,0,0,0,0,0,0,6,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,24,24,3,3,3,24,24,24,24,24,24,24,24,0,0,0},
'{0,0,0,0,0,0,0,24,24,24,24,24,24,24,24,24,24,24,24,24,24,0,0,0},
'{0,0,0,0,0,0,24,24,25,25,25,25,24,24,24,3,3,3,3,3,3,3,3,0},
'{0,0,0,0,0,24,24,25,25,25,3,24,24,24,25,24,25,24,25,24,0,0,0,0},
'{0,0,0,0,24,24,25,25,25,25,3,3,24,25,25,24,25,24,25,24,0,0,0,0},
'{0,0,0,0,0,24,24,25,25,25,3,24,24,24,25,24,25,24,25,24,0,0,0,0},
'{0,0,0,0,0,0,24,24,25,25,25,25,24,24,24,3,3,3,3,3,3,3,3,0},
'{0,0,0,0,0,0,0,24,24,24,24,24,24,24,24,24,24,24,24,24,24,0,0,0},
'{0,0,0,0,0,0,0,0,24,24,3,3,3,24,24,24,24,24,24,24,24,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,6,0,0,0,0,0,0,6,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,6,6,6,0,0,0,0,0,6,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,6,6,6,0,0,0,6,6,6,6,6,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,6,6,6,6,6,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};

	end
	
	always_ff
	begin
		data = carleft[DY][DX];
	//unique case (dir)
		//1'd0: data = truckleft[DY][DX];
		//1'd1: data = truckright[DY][DX];
		
	//endcase

	end
endmodule
