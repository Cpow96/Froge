module connrom
(
	input logic [5:0] DX, DY,
	output logic [7:0] data
);
// 1
	int conn [24][24];
	
	always_ff
	begin
	
	conn = '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0},
'{0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0},
'{0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0},
'{0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0},
'{0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0},
'{0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0},
'{0,0,0,0,1,1,29,1,1,1,1,1,1,1,1,1,29,1,1,1,0,0,0,0},
'{0,0,0,0,1,1,29,29,1,1,29,1,1,1,29,29,29,29,29,1,0,0,0,0},
'{0,0,0,0,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0},
'{0,0,0,0,29,29,29,5,5,5,29,29,29,29,5,5,5,29,29,29,0,0,0,0},
'{0,0,0,0,29,29,29,5,5,5,29,29,29,29,5,5,5,29,29,29,0,0,0,0},
'{0,0,0,0,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0},
'{0,0,0,0,29,29,29,29,6,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0},
'{0,0,0,0,29,29,29,29,6,6,29,29,29,6,6,29,29,29,29,29,0,0,0,0},
'{0,0,0,0,29,29,29,29,29,6,6,6,6,6,29,29,29,29,29,0,0,0,0,0},
'{0,0,0,0,0,29,29,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0},
'{0,0,0,0,0,0,29,29,29,29,29,29,29,29,29,29,29,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};

	end
	
	always_ff
	begin
		data = conn[DY][DX];
	//unique case (dir)
		//1'd0: data = truckleft[DY][DX];
		//1'd1: data = truckright[DY][DX];
		
	//endcase

	end
endmodule