module othercarrightrom
(
	input logic [5:0] DX, DY,
	input logic  dir,
	output logic [7:0] data
);
// 1
	int othercarright [24][32];
	
	always_ff
	begin
	
	othercarright = '{'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,23,23,23,23,0,0,0,0,0,0,0,0,0,0,0,0,0,0,23,23,23,23,0,0,0,0,0},
'{0,0,0,0,0,23,23,23,23,0,0,0,0,0,0,0,0,0,0,0,0,0,0,23,23,23,23,0,0,0,0,0},
'{0,0,0,0,21,23,23,23,23,21,21,21,0,0,0,0,0,0,0,20,20,21,21,23,23,23,23,21,21,0,0,0},
'{3,3,3,3,21,21,21,21,21,21,21,21,21,0,0,0,0,0,20,20,20,21,21,21,0,0,0,0,21,0,0,0},
'{0,0,3,3,20,20,20,20,20,20,21,21,21,21,21,20,20,20,20,3,20,21,21,21,0,0,21,21,21,21,0,0},
'{0,0,3,20,22,22,22,22,22,20,21,21,21,21,21,20,20,20,20,3,20,20,21,21,21,21,21,21,21,3,3,0},
'{0,0,3,20,22,22,22,22,22,20,21,21,21,21,21,20,19,20,20,20,20,20,20,25,25,25,25,25,25,3,3,0},
'{0,0,3,20,22,22,22,22,22,20,21,21,21,21,19,19,19,20,20,20,20,20,20,20,20,20,20,20,20,20,3,0},
'{0,0,3,20,22,22,22,22,22,20,21,21,21,21,19,19,19,20,20,20,20,20,19,19,19,19,19,19,19,20,3,0},
'{0,0,3,20,22,22,22,22,22,20,21,21,21,21,19,19,19,20,20,20,20,20,20,20,20,20,20,20,20,20,3,0},
'{0,0,3,20,22,22,22,22,22,20,21,21,21,21,21,20,19,20,20,20,20,20,20,25,25,25,25,25,25,3,3,0},
'{0,0,3,20,22,22,22,22,22,20,21,21,21,21,21,20,20,20,20,3,20,20,21,21,21,21,21,21,21,3,3,0},
'{0,0,3,3,20,20,20,20,20,20,21,21,21,21,21,20,20,20,20,3,20,21,21,21,0,0,21,21,21,21,0,0},
'{3,3,3,3,21,21,21,21,21,21,21,21,21,0,0,0,0,0,20,20,20,21,21,21,0,0,0,0,21,0,0,0},
'{0,0,0,0,21,23,23,23,23,21,21,21,0,0,0,0,0,0,0,20,20,21,21,23,23,23,23,21,21,0,0,0},
'{0,0,0,0,0,23,23,23,23,0,0,0,0,0,0,0,0,0,0,0,0,0,0,23,23,23,23,0,0,0,0,0},
'{0,0,0,0,0,23,23,23,23,0,0,0,0,0,0,0,0,0,0,0,0,0,0,23,23,23,23,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}};

	end
	
	always_ff
	begin
		data = othercarright[DY][DX];
	//unique case (dir)
		//1'd0: data = truckleft[DY][DX];
		//1'd1: data = truckright[DY][DX];
		
	//endcase

	end
endmodule