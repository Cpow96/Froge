module map_ROM_16
(
	input logic [9:0] currX, currY,
	output logic [7:0] outR, outG, outB
);
	// # of map sprites: 33 6'd
	// this array holds information on how the map is pieced together from sprites; numbers indicate different sprites of the map
	parameter bit [5:0] map_Layout [0:29][27:0] = '{'{6'd0, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd19, 6'd20, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd2},				// row 0
													 '{6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7},								// row 1
													 '{6'd3, 6'd4, 6'd8, 6'd9, 6'd9, 6'd10, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd5, 6'd6, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd8, 6'd9, 6'd9, 6'd10, 6'd4, 6'd7},							// row 2
													 '{6'd3, 6'd4, 6'd5, 6'd4, 6'd4, 6'd6, 6'd4, 6'd5, 6'd4, 6'd4, 6'd4, 6'd6, 6'd4, 6'd5, 6'd6, 6'd4, 6'd5, 6'd4, 6'd4, 6'd4, 6'd6, 6'd4, 6'd5, 6'd4, 6'd4, 6'd6, 6'd4, 6'd7},								// row 3
													 '{6'd3, 6'd4, 6'd11, 6'd12, 6'd12, 6'd13, 6'd4, 6'd11, 6'd12, 6'd12, 6'd12, 6'd13, 6'd4, 6'd11, 6'd13, 6'd4, 6'd11, 6'd12, 6'd12, 6'd12, 6'd13, 6'd4, 6'd11, 6'd12, 6'd12, 6'd13, 6'd4, 6'd7},		// row 4
													 '{6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7},								// row 5
													 '{6'd3, 6'd4, 6'd8, 6'd9, 6'd9, 6'd10, 6'd4, 6'd8, 6'd10, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd8, 6'd10, 6'd4, 6'd8, 6'd9, 6'd9, 6'd10, 6'd4, 6'd7},							// row 6
													 '{6'd3, 6'd4, 6'd11, 6'd12, 6'd12, 6'd13, 6'd4, 6'd5, 6'd6, 6'd4, 6'd11, 6'd12, 6'd12, 6'd21, 6'd22, 6'd12, 6'd12, 6'd13, 6'd4, 6'd5, 6'd6, 6'd4, 6'd11, 6'd12, 6'd12, 6'd13, 6'd4, 6'd7},			// row 7
													 '{6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7},								// row 8
													 '{6'd14, 6'd15, 6'd15, 6'd15, 6'd15, 6'd10, 6'd4, 6'd5, 6'd16, 6'd9, 6'd9, 6'd10, 6'd4, 6'd5, 6'd6, 6'd4, 6'd8, 6'd9, 6'd9, 6'd17, 6'd6, 6'd4, 6'd8, 6'd15, 6'd15, 6'd15, 6'd15, 6'd18},				// row 9
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd5, 6'd22, 6'd12, 6'd12, 6'd13, 6'd4, 6'd11, 6'd13, 6'd4, 6'd11, 6'd12, 6'd12, 6'd21, 6'd6, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},					// row 10
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},								// row 11
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd11, 6'd13, 6'd4, 6'd23, 6'd15, 6'd24, 6'd25, 6'd25, 6'd26, 6'd15, 6'd27, 6'd4, 6'd11, 6'd13, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},				// row 12
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},								// row 13
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd8, 6'd10, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd8, 6'd10, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},								// row 14
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd5, 6'd6, 6'd4, 6'd28, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd1, 6'd29, 6'd4, 6'd5, 6'd6, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},								// row 15
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},								// row 16
													 '{6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd3, 6'd4, 6'd5, 6'd6, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd5, 6'd6, 6'd4, 6'd7, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4},								// row 17
													 '{6'd0, 6'd1, 6'd1, 6'd1, 6'd1, 6'd13, 6'd4, 6'd11, 6'd13, 6'd4, 6'd11, 6'd12, 6'd12, 6'd21, 6'd22, 6'd12, 6'd12, 6'd13, 6'd4, 6'd11, 6'd13, 6'd4, 6'd11, 6'd1, 6'd1, 6'd1, 6'd1, 6'd2},				// row 18
													 '{6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7},								// row 19
													 '{6'd3, 6'd4, 6'd8, 6'd9, 6'd9, 6'd10, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd5, 6'd6, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd8, 6'd9, 6'd9, 6'd10, 6'd4, 6'd7},							// row 20
													 '{6'd3, 6'd4, 6'd11, 6'd12, 6'd21, 6'd6, 6'd4, 6'd11, 6'd12, 6'd12, 6'd12, 6'd13, 6'd4, 6'd11, 6'd13, 6'd4, 6'd11, 6'd12, 6'd12, 6'd12, 6'd13, 6'd4, 6'd5, 6'd22, 6'd12, 6'd13, 6'd4, 6'd7},		// row 21
													 '{6'd3, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd7},								// row 22
													 '{6'd30, 6'd9, 6'd10, 6'd4, 6'd5, 6'd6, 6'd4, 6'd8, 6'd10, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd8, 6'd10, 6'd4, 6'd5, 6'd6, 6'd4, 6'd8, 6'd9, 6'd31},						// row 23
													 '{6'd32, 6'd12, 6'd13, 6'd4, 6'd11, 6'd13, 6'd4, 6'd5, 6'd6, 6'd4, 6'd11, 6'd12, 6'd12, 6'd21, 6'd22, 6'd12, 6'd12, 6'd13, 6'd4, 6'd5, 6'd6, 6'd4, 6'd11, 6'd13, 6'd4, 6'd11, 6'd12, 6'd33},		// row 24
													 '{6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd5, 6'd6, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7},								// row 25
													 '{6'd3, 6'd4, 6'd8, 6'd9, 6'd9, 6'd9, 6'd9, 6'd17, 6'd16, 6'd9, 6'd9, 6'd10, 6'd4, 6'd5, 6'd6, 6'd4, 6'd8, 6'd9, 6'd9, 6'd17, 6'd16, 6'd9, 6'd9, 6'd9, 6'd9, 6'd10, 6'd4, 6'd7},						// row 26
													 '{6'd3, 6'd4, 6'd11, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd13, 6'd4, 6'd11, 6'd13, 6'd4, 6'd11, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd12, 6'd13, 6'd4, 6'd7},	// row 27
													 '{6'd3, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd4, 6'd7},								// row 28
													 '{6'd14, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd15, 6'd18}};	// row 29							// row 28
													 											 

	parameter [0:15][15:0] map_0 = {16'b0000000011111111,
											16'b0000000011111111,
											16'b0000111100000000,
											16'b0000111100000000,
											16'b0011000000000000,
											16'b0011000000000000,
											16'b0011000000111111,
											16'b0011000000111111,
											16'b1100000011000000,
											16'b1100000011000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000};
			
		
	parameter [0:15][15:0] map_1 = {16'b1111111111111111,
											16'b1111111111111111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
											

	parameter [0:15][15:0] map_19 = {16'b1111111111111111,
											 16'b1111111111111111,
											 16'b0000000000000000,
											 16'b0000000000000000,
											 16'b0000000000000000,
											 16'b0000000000000000,
											 16'b1111110000000000,
											 16'b1111110000000000,
											 16'b0000001100000000,
											 16'b0000001100000000,
											 16'b0000000011000000,
											 16'b0000000011000000,
											 16'b0000000011000000,
											 16'b0000000011000000,
											 16'b0000000011000000,
											 16'b0000000011000000};



	parameter [0:15][15:0] map_20 = {16'b1111111111111111,
											 16'b1111111111111111,
											 16'b0000000000000000,
											 16'b0000000000000000,
											 16'b0000000000000000,
											 16'b0000000000000000,
											 16'b0000000000111111,
											 16'b0000000000111111,
											 16'b0000000011000000,
											 16'b0000000011000000,
											 16'b0000001100000000,
											 16'b0000001100000000,
											 16'b0000001100000000,
											 16'b0000001100000000,
											 16'b0000001100000000,
											 16'b0000001100000000};
											 

	parameter [0:15][15:0] map_2 = {16'b1111111100000000,
											16'b1111111100000000,
											16'b0000000011110000,
											16'b0000000011110000,
											16'b0000000000001100,
											16'b0000000000001100,
											16'b1111110000001100,
											16'b1111110000001100,
											16'b0000001100000011,
											16'b0000001100000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,	
											16'b0000000011000011};
										

	parameter [0:15][15:0] map_4 = {16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111};
		
	parameter [0:15][15:0] map_3 = {16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000};
										
	parameter [0:15][15:0] map_5 = {16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000};

	parameter [0:15][15:0] map_6 = {16'b0000001100000000,		
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000,	
											16'b0000001100000000};
										
	parameter [0:15][15:0] map_7 = {16'b0000000011000011,		
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011};
									
	parameter [0:15][15:0] map_8 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000001111,
											16'b0000000000001111,
											16'b0000000000110000,
											16'b0000000000110000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000};
									
	parameter [0:15][15:0] map_9 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
									
	parameter [0:15][15:0] map_10 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111000000000000,
											16'b1111000000000000,
											16'b0000110000000000,
											16'b0000110000000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											};
							
	parameter [0:15][15:0] map_11 = {16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000000110000,
											16'b0000000000110000,
											16'b0000000000001111,
											16'b0000000000001111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
						
	parameter [0:15][15:0] map_12 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
					
	parameter [0:15][15:0] map_13 = {16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000110000000000,
											16'b0000110000000000,
											16'b1111000000000000,
											16'b1111000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
											
	parameter [0:15][15:0] map_21 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111110000000000,
											16'b1111110000000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000};
											
	parameter [0:15][15:0] map_22 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000111111,
											16'b0000000000111111,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000};
											
	parameter [0:15][15:0] map_14 = {16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100000011000000,
											16'b1100000011000000,
											16'b0011000000111111,
											16'b0011000000111111,
											16'b0011000000000000,
											16'b0011000000000000,
											16'b0000111100000000,
											16'b0000111100000000,
											16'b0000000011111111,
											16'b0000000011111111};
											
	parameter [0:15][15:0] map_15 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111};
											
	parameter [0:15][15:0] map_16 = {16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000000111111,
											16'b0000000000111111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
											
	parameter [0:15][15:0] map_17 = {16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b1111110000000000,
											16'b1111110000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
											
	parameter [0:15][15:0] map_18 = {16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000001100000011,
											16'b0000001100000011,
											16'b1111110000001100,
											16'b1111110000001100,
											16'b0000000000001100,
											16'b0000000000001100,
											16'b0000000011110000,
											16'b0000000011110000,
											16'b1111111100000000,
											16'b1111111100000000};

	parameter [0:15][15:0] map_23 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000011111111,
											16'b0000000011111111,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000011,
											16'b0000000011000011};
											
	parameter [0:15][15:0] map_24 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b1111111111111111,
											16'b1111111111111111};
											
	parameter [0:15][15:0] map_25 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b0000000000000000,
											16'b0000000000000000};
											
	parameter [0:15][15:0] map_26 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111111111111,
											16'b1111111111111111,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1111111111111111,
											16'b1111111111111111};
											
	parameter [0:15][15:0] map_27 = {16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b1111111100000000,
											16'b1111111100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b1100001100000000,
											16'b1100001100000000};

	parameter [0:15][15:0] map_28 = {16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011000000,
											16'b0000000011111111,
											16'b0000000011111111,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
											
	parameter [0:15][15:0] map_29 = {16'b1100001100000000,
											16'b1100001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b0000001100000000,
											16'b1111111100000000,
											16'b1111111100000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000,
											16'b0000000000000000};
											
	parameter [0:15][15:0] map_30 = {16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100000011000000,
											16'b1100000011000000,
											16'b1100000000111111,
											16'b1100000000111111,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000};
											
	parameter [0:15][15:0] map_31 = {16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000001100000011,
											16'b0000001100000011,
											16'b1111110000000011,
											16'b1111110000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011};

	parameter [0:15][15:0] map_32 = {16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000000000,
											16'b1100000000111111,
											16'b1100000000111111,
											16'b1100000011000000,
											16'b1100000011000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000,
											16'b1100001100000000};
											
	parameter [0:15][15:0] map_33 = {16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b0000000000000011,
											16'b1111110000000011,
											16'b1111110000000011,
											16'b0000001100000011,
											16'b0000001100000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011,
											16'b0000000011000011};
											
// 1
//	assign data = mapROM[addr];

	// translate coordinates to a 40x30 grid system
	logic [15:0] indexX, indexY;
	logic [5:0] mapSprite;
	logic [9:0] x, y;
	logic [15:0] spriteData;
	assign y = currY >> 10'd4;
	assign x = currX >> 10'd4;
	assign indexX = {6'b0, currX & 10'd15};//currX % 10'd8;
	assign indexY = {6'b0, currY & 10'd15};//currY % 10'd8;
//	assign indexX = currX % 10'd8;
//	assign indexY = currY % 10'd8;
	assign mapSprite = map_Layout[y][27-x];
//   assign mapSprite = 6'd1;
	
	always_comb begin
	spriteData = 8'd0;
	unique case (mapSprite)
		6'd0: begin
			spriteData = map_0[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd1: begin
			spriteData = map_1[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd2: begin
			spriteData = map_2[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd19: begin
			spriteData = map_19[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd20: begin
			spriteData = map_20[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd3: begin
			spriteData = map_3[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end	
		
		6'd4: begin
			spriteData = map_4[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd5: begin
			spriteData = map_5[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd6: begin
			spriteData = map_6[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd7: begin
			spriteData = map_7[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd8: begin
			spriteData = map_8[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd9: begin
			spriteData = map_9[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd10: begin
			spriteData = map_10[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd11: begin
			spriteData = map_11[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd12: begin
			spriteData = map_12[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd13: begin
			spriteData = map_13[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
	
		6'd21: begin
			spriteData = map_21[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd22: begin
			spriteData = map_22[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end			

		6'd14: begin
			spriteData = map_14[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd15: begin
			spriteData = map_15[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd16: begin
			spriteData = map_16[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd17: begin
			spriteData = map_17[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd18: begin
			spriteData = map_18[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd23: begin
			spriteData = map_23[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd24: begin
			spriteData = map_24[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd25: begin
			spriteData = map_25[indexY];
			if (spriteData[15-indexX])
			begin
				// pink
				outR = 8'hff;
				outG = 8'hc0;
				outB = 8'hcb;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd26: begin
			spriteData = map_26[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd27: begin
			spriteData = map_27[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end
		
		6'd28: begin
			spriteData = map_28[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end

		6'd29: begin
			spriteData = map_29[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end	

		6'd30: begin
			spriteData = map_30[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end		

		6'd31: begin
			spriteData = map_31[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end	
		
		6'd32: begin
			spriteData = map_32[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end	

		6'd33: begin
			spriteData = map_33[indexY];
			if (spriteData[15-indexX])
			begin
				// blue
				outR = 8'h00;
				outG = 8'h00;
				outB = 8'hff;
			end
			else
			begin
				outR = 8'h3f;
				outG = 8'h00;
				outB = 8'h3f;
			end
		end	
		
		default: begin
			outR = 8'hff;
			outG = 8'hff;
			outB = 8'hff;
		end
	endcase
	end
	
endmodule